module filtrosvga(
	input logic clk, rst,
	input logic [7:0] datain,
	output logic [7:0] dataout
);

